-- ----------------------------------------------------------------------------
-- Author     : Michael Jørgensen
-- Platform   : AMD Artix 7
-- ----------------------------------------------------------------------------
-- Description:
-- ----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package wbus_pkg is

  type slv32_array_type is array (natural range <>) of std_logic_vector(31 downto 0);

end package wbus_pkg;

package body wbus_pkg is

end package body wbus_pkg;

