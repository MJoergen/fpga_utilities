-- ---------------------------------------------------------------------------------------
-- Description:
-- ---------------------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package axip_pkg is

  subtype nat16_type is natural range 0 to 65535;

  type nat16_array_type is array (natural range <>) of nat16_type;

end package axip_pkg;


package body axip_pkg is

end package body axip_pkg;

